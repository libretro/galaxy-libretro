BSV1    s��    